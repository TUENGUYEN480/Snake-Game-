module top (
  input logic clk_i,
    input logic reset_i,
	 input logic enter_i,
    input logic KEY_0, KEY_1, KEY_2, KEY_3,
	 output logic [6:0] hang_chuc,
	 output logic [6:0] hang_don_vi,
    output logic hsync,
    output logic vsync,
    output logic display_on,
    output logic vga_clk,
    output logic [7:0] r_o,
    output logic [7:0] g_o,
    output logic [7:0] b_o
);
	 logic update_clk;
    logic [3:0] direction;
    logic [9:0] hpos, vpos;
    logic head_snake_gfx, body_snake_gfx, apple_gfx, border_gfx;
    logic snake_colline, playing,enter, game_over,apple_colline_o;

   key_board key_inst (
        .clk_i(clk_i),
		  .reset(reset_i),
        .KEY_0(KEY_0),
        .KEY_1(KEY_1),
        .KEY_2(KEY_2),
        .KEY_3(KEY_3),
        .direction_o(direction)
    );
    //module clk_VGA
	 clk_VGA clk_VGA1(
	     .clk_i(clk_i),
		  .clk_vga(vga_clk)
	 );
    // Module speed_control
    speed_control speed_inst (
        .clk_i(clk_i),
        
        .update_clk_o(update_clk)
    );

    // Module VGA_controller
    VGA_controller vga_inst (
        .clk_i(vga_clk),
        .reset(reset_i),
        .hsync(hsync),
        .vsync(vsync),
        .display_on_o(display_on),
        .hpos(hpos),
        .vpos(vpos)
    );

    // Module game_state_machine
    game_stage_machine state_inst (
        .clk_i(vga_clk),
        .reset_i(reset_i),
        .snake_colline_i(snake_colline),
        .enter_i(enter_i),
        .playing_o(playing),
        .game_over_o(game_over)
    );

    // Module snake_and_apple
    snake_and_apple snake_inst (
        .clk_i(vga_clk),
        .snake_clk_i(update_clk),
        .reset_i(reset_i),
        .direction_i(direction),
		  .enter_i(enter_i),
        .hpos_i(hpos),
        .vpos_i(vpos),
        .playing_i(playing),
        .game_over_i(game_over),
        .snake_colline_o(snake_colline),
		  .apple_colline_o (apple_colline_o),
        .head_snake_gfx_o(head_snake_gfx),
        .body_snake_gfx_o(body_snake_gfx),
        .apple_gfx_o(apple_gfx),
        .border_gfx_o(border_gfx)
    );

    // Module drawer
    drawer draw_inst (
        .display_enable_i(display_on),
        .head_snake_gfx_i(head_snake_gfx),
        .body_snake_gfx_i(body_snake_gfx),
        .apple_gfx_i(apple_gfx),
        .border_gfx_i(border_gfx),
        .r_o(r_o),
        .g_o(g_o),
        .b_o(b_o)
    );

	 led_7_doan led_7_doan_inst (
		.clk_i(clk_i),      
      .reset_i(reset_i),   
   	.apple_colline(apple_colline_o), 
      .hang_chuc(hang_chuc), 
      .hang_don_vi(hang_don_vi),
	);
endmodule
	